library verilog;
use verilog.vl_types.all;
entity counter is
end counter;
