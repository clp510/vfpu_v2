library verilog;
use verilog.vl_types.all;
entity vfpu_dc_pkg is
end vfpu_dc_pkg;
