library verilog;
use verilog.vl_types.all;
entity top_tb_m is
end top_tb_m;
