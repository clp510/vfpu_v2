library verilog;
use verilog.vl_types.all;
entity test_dutw_if is
    port(
        clk             : in     vl_logic
    );
end test_dutw_if;
