library verilog;
use verilog.vl_types.all;
entity top_tb_m_sv_unit is
end top_tb_m_sv_unit;
