library verilog;
use verilog.vl_types.all;
entity mul_24x24_tb is
end mul_24x24_tb;
