//==================================================================
//File Name	: vfpu_top_m.sv
//Author	: clp
//Email		: clp510@tju.edu.cn
//Date		: 2015.01.09
//Revision	: v1.0
//Description: top level module of vfpu verification platform
// 1) instance DUT module and SV program
// 2) generate clk and rst_n signal
//------------------------------------------------------------
//Copyright(c)by VLSI lab of Tianjin university
//all rights reserved
//==================================================================

`timescale 1ns/1ns
//`define MAX_NUM 1000

import vfpu_dc_pkg::BIT ;

module  top_tb_m();


BIT         clk;
BIT         rst_n;

//interface between DUT and SV platform
test_dutw_if    test_dutw_if_inst( clk );

//generate clk and rst_n signal
initial
begin
    clk     = 1'b1;
    forever #5 clk = ~clk;
end


//connect the clock signal
//assign  test_dutw_if_inst.clk  = clk;
/*
initial
begin
    $monitor($time,"test_dutw_if_inst.clk=%b\n",clk);
end   
*/ 
//reset signal should be generated by test program
//--------------------------------------------------
//instance test program
test_p    test_p_inst   (
                    clk,
                   test_dutw_if_inst
                   );
//instance dut_wrapper module
dut_wrapper_m dut_wrapper_m_inst    (
                                clk,
                                test_dutw_if_inst
                                );
endmodule                               

