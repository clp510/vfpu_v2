library verilog;
use verilog.vl_types.all;
entity dut_wrapper_m_sv_unit is
end dut_wrapper_m_sv_unit;
