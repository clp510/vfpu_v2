library verilog;
use verilog.vl_types.all;
entity test_p_sv_unit is
end test_p_sv_unit;
