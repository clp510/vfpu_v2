library verilog;
use verilog.vl_types.all;
entity dut_wrapper_m is
    port(
        clk             : in     vl_logic
    );
end dut_wrapper_m;
