library verilog;
use verilog.vl_types.all;
entity maf_tb is
end maf_tb;
