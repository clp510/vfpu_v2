library verilog;
use verilog.vl_types.all;
entity vfpu_if_sv_unit is
end vfpu_if_sv_unit;
