library verilog;
use verilog.vl_types.all;
entity test_p is
    port(
        clk             : in     vl_logic
    );
end test_p;
